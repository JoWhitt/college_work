INFO:HDLCompiler:1061 - Parsing VHDL file "U:/Comp_Arch/Register.vhd" into library work
ERROR:HDLCompiler:806 - "U:/Comp_Arch/Register.vhd" Line 32: Syntax error near "register".
ERROR:HDLCompiler:806 - "U:/Comp_Arch/Register.vhd" Line 39: Syntax error near "register".
INFO:HDLCompiler:1061 - Parsing VHDL file "U:/Comp_Arch/decoder_2to4.vhd" into library work
ERROR:HDLCompiler:806 - "U:/Comp_Arch/decoder_2to4.vhd" Line 36: Syntax error near "end".
INFO:HDLCompiler:1061 - Parsing VHDL file "U:/Comp_Arch/mux2_4bit.vhd" into library work
ERROR:HDLCompiler:806 - "U:/Comp_Arch/mux2_4bit.vhd" Line 40: Syntax error near "Z".
ERROR:ProjectMgmt - 4 error(s) found while parsing design hierarchy.
